module RCA4 (input  logic[3:0] a, b, input logic cin, output logic cout, sum);
   output logic cout[1], cout[2], cout[3];
   
  
   
endmodule
